--//////////////////////////////////////////////////////////////////////////////
-- Project Name:	CoCo3FPGA Version 4.0
-- File Name:		CoCo_ram_128x8.vhd
--
-- CoCo3 in an FPGA
--
-- Revision: 5.x.x
--//////////////////////////////////////////////////////////////////////////////
--
-- Color Computer 3 compatible system on a chip
--
-- Version : 5.0.x.x
--
-- Copyright (c) 2008 Gary Becker (gary_l_becker@yahoo.com)
--
-- All rights reserved
--
-- Redistribution and use in source and synthezised forms, with or without
-- modification, are permitted provided that the following conditions are met:
--
-- Redistributions of source code must retain the above copyright notice,
-- this list of conditions and the following disclaimer.
--
-- Redistributions in synthesized form must reproduce the above copyright
-- notice, this list of conditions and the following disclaimer in the
-- documentation and/or other materials provided with the distribution.
--
-- Neither the name of the author nor the names of other contributors may
-- be used to endorse or promote products derived from this software without
-- specific prior written permission.
--
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
-- AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR
-- PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE AUTHOR OR CONTRIBUTORS BE
-- LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
-- CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
-- SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
-- INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
-- CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
-- POSSIBILITY OF SUCH DAMAGE.
--
-- Please report bugs to the author, but before you do so, please
-- make sure that this is not a derivative work and that
-- you have the latest version of this file.
--
-- The latest version of this file can be found at:
--      http://groups.yahoo.com/group/CoCo3FPGA
--
-- File history :
--
--  1.0			Full Release
--  2.0			Partial Release
--  3.0			Full Release
--  3.0.0.1		Update to fix DoD interrupt issue
--//////////////////////////////////////////////////////////////////////////////
-- Gary Becker
-- gary_L_becker@yahoo.com
--//////////////////////////////////////////////////////////////////////////////
--//////////////////////////////////////////////////////////////////////////////
--////////////////////////////////////////////////////////////////////////////////
--// MISTer Conversion by Stan Hodge and Alan Steremberg (& Gary Becker)
--// stan.pda@gmail.com
--// 
--////////////////////////////////////////////////////////////////////////////////


library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

entity COCO_SRAM_6116 is
  port (
	CLK				: in	std_logic;
	ENA				: in 	std_logic;
    ADDR        	: in    std_logic_vector(6 downto 0);
	R_W				: in	std_logic;
	DATA_I			: in	std_logic_vector(7 downto 0);
    DATA_O        	: out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of COCO_SRAM_128x8 is

  type SRAM_ARRAY is array(0 to 127) of std_logic_vector(7 downto 0);
  signal SRAM : SRAM_ARRAY;

begin

  P_SRAM : process(CLK,ADDR,R_W,DATA_I)
  begin
	if CLK'event and CLK='1' then
		if ENA = '1' and R_W = '0' then
    		SRAM(to_integer(unsigned(ADDR))) <= DATA_I;
		end if;
	end if;
  end process;

  DATA_O <= SRAM(to_integer(unsigned(ADDR)));

end RTL;
