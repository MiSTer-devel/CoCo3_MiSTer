-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

entity coco3_Char_ROM is
  port (
    RD_CLK      : in    std_logic;
    ADDR_R      : in    std_logic_vector(11 downto 0);
    DATA_R      : out   std_logic_vector(7 downto 0);

    WR_CLK      : in    std_logic;
	WE			: in    std_logic;
    ADDR_W      : in    std_logic_vector(11 downto 0);
    DATA_W      : in    std_logic_vector(7 downto 0)
    );
end;

architecture RTL of coco3_Char_ROM is


  type RAM_ARRAY is array(0 to 4095) of std_logic_vector(7 downto 0);
  signal RAM : RAM_ARRAY := (
    x"1C",x"22",x"20",x"20",x"20",x"22",x"1C",x"08", -- 0x0000
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0008
    x"22",x"00",x"22",x"22",x"22",x"26",x"1A",x"00", -- 0x0010
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0018
    x"04",x"08",x"1C",x"22",x"3E",x"20",x"1C",x"00", -- 0x0020
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0028
    x"08",x"14",x"1C",x"02",x"1E",x"22",x"1E",x"00", -- 0x0030
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0038
    x"14",x"00",x"1C",x"02",x"1E",x"22",x"1E",x"00", -- 0x0040
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0048
    x"10",x"08",x"1C",x"02",x"1E",x"22",x"1E",x"00", -- 0x0050
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0058
    x"08",x"00",x"1C",x"02",x"1E",x"22",x"1E",x"00", -- 0x0060
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0068
    x"00",x"00",x"1C",x"22",x"20",x"22",x"1C",x"08", -- 0x0070
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0078
    x"08",x"14",x"1C",x"22",x"3E",x"20",x"1C",x"00", -- 0x0080
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0088
    x"14",x"00",x"1C",x"22",x"3E",x"20",x"1C",x"00", -- 0x0090
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0098
    x"10",x"08",x"1C",x"22",x"3E",x"20",x"1C",x"00", -- 0x00A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00A8
    x"14",x"00",x"18",x"08",x"08",x"08",x"1C",x"00", -- 0x00B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00B8
    x"08",x"14",x"00",x"18",x"08",x"08",x"1C",x"00", -- 0x00C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00C8
    x"00",x"0C",x"12",x"1C",x"12",x"12",x"1C",x"20", -- 0x00D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00D8
    x"22",x"08",x"14",x"22",x"3E",x"22",x"22",x"00", -- 0x00E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00E8
    x"08",x"08",x"14",x"22",x"3E",x"22",x"22",x"00", -- 0x00F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00F8
    x"04",x"08",x"1C",x"22",x"22",x"22",x"1C",x"00", -- 0x0100
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0108
    x"00",x"00",x"34",x"0A",x"1E",x"28",x"1E",x"00", -- 0x0110
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0118
    x"1E",x"28",x"28",x"3C",x"28",x"28",x"2C",x"00", -- 0x0120
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0128
    x"08",x"14",x"1C",x"22",x"22",x"22",x"1C",x"00", -- 0x0130
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0138
    x"14",x"00",x"1C",x"22",x"22",x"22",x"1C",x"00", -- 0x0140
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0148
    x"00",x"00",x"1C",x"26",x"2E",x"32",x"1C",x"00", -- 0x0150
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0158
    x"08",x"14",x"00",x"22",x"22",x"26",x"1A",x"00", -- 0x0160
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0168
    x"10",x"08",x"22",x"22",x"22",x"26",x"1A",x"00", -- 0x0170
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0178
    x"1C",x"26",x"2A",x"2A",x"2A",x"32",x"1C",x"00", -- 0x0180
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0188
    x"22",x"1C",x"22",x"22",x"22",x"22",x"1C",x"00", -- 0x0190
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0198
    x"14",x"22",x"22",x"22",x"22",x"22",x"1C",x"00", -- 0x01A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01A8
    x"1C",x"20",x"1C",x"22",x"1C",x"02",x"1C",x"00", -- 0x01B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01B8
    x"04",x"0A",x"08",x"1C",x"08",x"0A",x"3C",x"00", -- 0x01C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01C8
    x"08",x"08",x"3E",x"08",x"08",x"00",x"3E",x"00", -- 0x01D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01D8
    x"04",x"0A",x"04",x"00",x"00",x"00",x"00",x"00", -- 0x01E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01E8
    x"04",x"0A",x"08",x"1C",x"08",x"08",x"28",x"10", -- 0x01F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0200
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0208
    x"08",x"08",x"08",x"08",x"08",x"00",x"08",x"00", -- 0x0210
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0218
    x"14",x"14",x"14",x"00",x"00",x"00",x"00",x"00", -- 0x0220
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0228
    x"14",x"14",x"3E",x"14",x"3E",x"14",x"14",x"00", -- 0x0230
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0238
    x"08",x"1E",x"28",x"1C",x"0A",x"3C",x"08",x"00", -- 0x0240
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0248
    x"32",x"32",x"04",x"08",x"10",x"26",x"26",x"00", -- 0x0250
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0258
    x"10",x"28",x"28",x"10",x"2A",x"24",x"1A",x"00", -- 0x0260
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0268
    x"08",x"08",x"10",x"00",x"00",x"00",x"00",x"00", -- 0x0270
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0278
    x"08",x"10",x"20",x"20",x"20",x"10",x"08",x"00", -- 0x0280
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0288
    x"08",x"04",x"02",x"02",x"02",x"04",x"08",x"00", -- 0x0290
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0298
    x"00",x"08",x"2A",x"1C",x"1C",x"2A",x"08",x"00", -- 0x02A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02A8
    x"00",x"08",x"08",x"3E",x"08",x"08",x"00",x"00", -- 0x02B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02B8
    x"00",x"00",x"00",x"00",x"00",x"08",x"08",x"10", -- 0x02C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02C8
    x"00",x"00",x"00",x"3E",x"00",x"00",x"00",x"00", -- 0x02D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"00", -- 0x02E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02E8
    x"00",x"02",x"04",x"08",x"10",x"20",x"00",x"00", -- 0x02F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02F8
    x"1C",x"22",x"26",x"2A",x"32",x"22",x"1C",x"00", -- 0x0300
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0308
    x"08",x"18",x"08",x"08",x"08",x"08",x"1C",x"00", -- 0x0310
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0318
    x"1C",x"22",x"02",x"1C",x"20",x"20",x"3E",x"00", -- 0x0320
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0328
    x"1C",x"22",x"02",x"04",x"02",x"22",x"1C",x"00", -- 0x0330
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0338
    x"04",x"0C",x"14",x"24",x"3E",x"04",x"04",x"00", -- 0x0340
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0348
    x"3E",x"20",x"3C",x"02",x"02",x"02",x"3C",x"00", -- 0x0350
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0358
    x"1C",x"20",x"20",x"3C",x"22",x"22",x"1C",x"00", -- 0x0360
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0368
    x"3E",x"02",x"04",x"08",x"10",x"20",x"20",x"00", -- 0x0370
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0378
    x"1C",x"22",x"22",x"1C",x"22",x"22",x"1C",x"00", -- 0x0380
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0388
    x"1C",x"22",x"22",x"1E",x"02",x"02",x"1C",x"00", -- 0x0390
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0398
    x"00",x"00",x"08",x"00",x"00",x"08",x"00",x"00", -- 0x03A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03A8
    x"00",x"00",x"08",x"00",x"00",x"08",x"08",x"10", -- 0x03B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03B8
    x"04",x"08",x"10",x"20",x"10",x"08",x"04",x"00", -- 0x03C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03C8
    x"00",x"00",x"3E",x"00",x"3E",x"00",x"00",x"00", -- 0x03D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03D8
    x"10",x"08",x"04",x"02",x"04",x"08",x"10",x"00", -- 0x03E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03E8
    x"1C",x"22",x"02",x"04",x"08",x"00",x"08",x"00", -- 0x03F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03F8
    x"1C",x"22",x"02",x"1A",x"2A",x"2A",x"1C",x"00", -- 0x0400
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0408
    x"08",x"14",x"22",x"22",x"3E",x"22",x"22",x"00", -- 0x0410
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0418
    x"3C",x"12",x"12",x"1C",x"12",x"12",x"3C",x"00", -- 0x0420
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0428
    x"1C",x"22",x"20",x"20",x"20",x"22",x"1C",x"00", -- 0x0430
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0438
    x"3C",x"12",x"12",x"12",x"12",x"12",x"3C",x"00", -- 0x0440
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0448
    x"3E",x"20",x"20",x"3C",x"20",x"20",x"3E",x"00", -- 0x0450
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0458
    x"3E",x"20",x"20",x"3C",x"20",x"20",x"20",x"00", -- 0x0460
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0468
    x"1E",x"20",x"20",x"26",x"22",x"22",x"1C",x"00", -- 0x0470
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0478
    x"22",x"22",x"22",x"3E",x"22",x"22",x"22",x"00", -- 0x0480
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0488
    x"1C",x"08",x"08",x"08",x"08",x"08",x"1C",x"00", -- 0x0490
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0498
    x"02",x"02",x"02",x"02",x"22",x"22",x"1C",x"00", -- 0x04A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04A8
    x"22",x"24",x"28",x"30",x"28",x"24",x"22",x"00", -- 0x04B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04B8
    x"20",x"20",x"20",x"20",x"20",x"20",x"3E",x"00", -- 0x04C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04C8
    x"22",x"36",x"2A",x"2A",x"22",x"22",x"22",x"00", -- 0x04D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04D8
    x"22",x"32",x"2A",x"26",x"22",x"22",x"22",x"00", -- 0x04E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04E8
    x"1C",x"22",x"22",x"22",x"22",x"22",x"1C",x"00", -- 0x04F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04F8
    x"3C",x"22",x"22",x"3C",x"20",x"20",x"20",x"00", -- 0x0500
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0508
    x"1C",x"22",x"22",x"22",x"2A",x"24",x"1A",x"00", -- 0x0510
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0518
    x"3C",x"22",x"22",x"3C",x"28",x"24",x"22",x"00", -- 0x0520
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0528
    x"1C",x"22",x"10",x"08",x"04",x"22",x"1C",x"00", -- 0x0530
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0538
    x"3E",x"08",x"08",x"08",x"08",x"08",x"08",x"00", -- 0x0540
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0548
    x"22",x"22",x"22",x"22",x"22",x"22",x"1C",x"00", -- 0x0550
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0558
    x"22",x"22",x"22",x"14",x"14",x"08",x"08",x"00", -- 0x0560
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0568
    x"22",x"22",x"22",x"2A",x"2A",x"36",x"22",x"00", -- 0x0570
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0578
    x"22",x"22",x"14",x"08",x"14",x"22",x"22",x"00", -- 0x0580
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0588
    x"22",x"22",x"14",x"08",x"08",x"08",x"08",x"00", -- 0x0590
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0598
    x"3E",x"02",x"04",x"08",x"10",x"20",x"3E",x"00", -- 0x05A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05A8
    x"38",x"20",x"20",x"20",x"20",x"20",x"38",x"00", -- 0x05B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05B8
    x"20",x"20",x"10",x"08",x"04",x"02",x"02",x"00", -- 0x05C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05C8
    x"0E",x"02",x"02",x"02",x"02",x"02",x"0E",x"00", -- 0x05D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05D8
    x"08",x"1C",x"2A",x"08",x"08",x"08",x"08",x"00", -- 0x05E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05E8
    x"00",x"08",x"10",x"3E",x"10",x"08",x"00",x"00", -- 0x05F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05F8
    x"08",x"14",x"22",x"00",x"00",x"00",x"00",x"00", -- 0x0600
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0608
    x"00",x"00",x"1C",x"02",x"1E",x"22",x"1E",x"00", -- 0x0610
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0618
    x"20",x"20",x"2C",x"32",x"22",x"32",x"2C",x"00", -- 0x0620
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0628
    x"00",x"00",x"1C",x"22",x"20",x"22",x"1C",x"00", -- 0x0630
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0638
    x"02",x"02",x"1A",x"26",x"22",x"26",x"1A",x"00", -- 0x0640
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0648
    x"00",x"00",x"1C",x"22",x"3E",x"20",x"1C",x"00", -- 0x0650
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0658
    x"04",x"0A",x"08",x"1C",x"08",x"08",x"08",x"00", -- 0x0660
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0668
    x"00",x"00",x"1A",x"26",x"26",x"1A",x"02",x"1C", -- 0x0670
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0678
    x"20",x"20",x"2C",x"32",x"22",x"22",x"22",x"00", -- 0x0680
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0688
    x"00",x"08",x"00",x"18",x"08",x"08",x"1C",x"00", -- 0x0690
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0698
    x"00",x"02",x"00",x"02",x"02",x"02",x"22",x"1C", -- 0x06A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06A8
    x"20",x"20",x"24",x"28",x"30",x"28",x"24",x"00", -- 0x06B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06B8
    x"18",x"08",x"08",x"08",x"08",x"08",x"1C",x"00", -- 0x06C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06C8
    x"00",x"00",x"14",x"2A",x"2A",x"2A",x"2A",x"00", -- 0x06D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06D8
    x"00",x"00",x"2C",x"32",x"22",x"22",x"22",x"00", -- 0x06E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06E8
    x"00",x"00",x"1C",x"22",x"22",x"22",x"1C",x"00", -- 0x06F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06F8
    x"00",x"00",x"2C",x"32",x"32",x"2C",x"20",x"20", -- 0x0700
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0708
    x"00",x"00",x"1A",x"26",x"26",x"1A",x"02",x"02", -- 0x0710
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0718
    x"00",x"00",x"2C",x"32",x"20",x"20",x"20",x"00", -- 0x0720
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0728
    x"00",x"00",x"1E",x"20",x"1C",x"02",x"3C",x"00", -- 0x0730
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0738
    x"10",x"10",x"38",x"10",x"10",x"12",x"0C",x"00", -- 0x0740
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0748
    x"00",x"00",x"22",x"22",x"22",x"26",x"1A",x"00", -- 0x0750
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0758
    x"00",x"00",x"22",x"22",x"22",x"14",x"08",x"00", -- 0x0760
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0768
    x"00",x"00",x"22",x"2A",x"2A",x"14",x"14",x"00", -- 0x0770
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0778
    x"00",x"00",x"22",x"14",x"08",x"14",x"22",x"00", -- 0x0780
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0788
    x"00",x"00",x"22",x"22",x"22",x"1E",x"02",x"1C", -- 0x0790
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0798
    x"00",x"00",x"3E",x"04",x"08",x"10",x"3E",x"00", -- 0x07A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07A8
    x"08",x"10",x"10",x"20",x"10",x"10",x"08",x"00", -- 0x07B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07B8
    x"08",x"08",x"08",x"00",x"08",x"08",x"08",x"00", -- 0x07C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07C8
    x"08",x"04",x"04",x"02",x"04",x"04",x"08",x"00", -- 0x07D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07D8
    x"10",x"2A",x"04",x"00",x"00",x"00",x"00",x"00", -- 0x07E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"3E",x"00", -- 0x07F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07F8
    x"00",x"00",x"1C",x"22",x"20",x"20",x"20",x"22", -- 0x0800
    x"1C",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0808
    x"00",x"00",x"22",x"00",x"22",x"22",x"22",x"26", -- 0x0810
    x"1A",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0818
    x"00",x"00",x"04",x"08",x"1C",x"22",x"3E",x"20", -- 0x0820
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0828
    x"00",x"00",x"08",x"14",x"1C",x"02",x"1E",x"22", -- 0x0830
    x"1E",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0838
    x"00",x"00",x"14",x"00",x"1C",x"02",x"1E",x"22", -- 0x0840
    x"1E",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0848
    x"00",x"00",x"10",x"08",x"1C",x"02",x"1E",x"22", -- 0x0850
    x"1E",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0858
    x"00",x"00",x"08",x"00",x"1C",x"02",x"1E",x"22", -- 0x0860
    x"1E",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0868
    x"00",x"00",x"00",x"00",x"1C",x"22",x"20",x"22", -- 0x0870
    x"1C",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0878
    x"00",x"00",x"08",x"14",x"1C",x"22",x"3E",x"20", -- 0x0880
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0888
    x"00",x"00",x"14",x"00",x"1C",x"22",x"3E",x"20", -- 0x0890
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0898
    x"00",x"00",x"10",x"08",x"1C",x"22",x"3E",x"20", -- 0x08A0
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x08A8
    x"00",x"00",x"14",x"00",x"18",x"08",x"08",x"08", -- 0x08B0
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x08B8
    x"00",x"00",x"08",x"14",x"00",x"18",x"08",x"08", -- 0x08C0
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x08C8
    x"00",x"00",x"00",x"0C",x"12",x"1C",x"12",x"12", -- 0x08D0
    x"1C",x"20",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x08D8
    x"00",x"00",x"22",x"08",x"14",x"22",x"3E",x"22", -- 0x08E0
    x"22",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x08E8
    x"00",x"00",x"08",x"08",x"14",x"22",x"3E",x"22", -- 0x08F0
    x"22",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x08F8
    x"00",x"00",x"04",x"08",x"1C",x"22",x"22",x"22", -- 0x0900
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0908
    x"00",x"00",x"00",x"00",x"34",x"0A",x"1E",x"28", -- 0x0910
    x"1E",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0918
    x"00",x"00",x"1E",x"28",x"28",x"3C",x"28",x"28", -- 0x0920
    x"2C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0928
    x"00",x"00",x"08",x"14",x"1C",x"22",x"22",x"22", -- 0x0930
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0938
    x"00",x"00",x"14",x"00",x"1C",x"22",x"22",x"22", -- 0x0940
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0948
    x"00",x"00",x"00",x"00",x"1C",x"26",x"2E",x"32", -- 0x0950
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0958
    x"00",x"00",x"08",x"14",x"00",x"22",x"22",x"26", -- 0x0960
    x"1A",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0968
    x"00",x"00",x"10",x"08",x"22",x"22",x"22",x"26", -- 0x0970
    x"1A",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0978
    x"00",x"00",x"1C",x"26",x"2A",x"2A",x"2A",x"32", -- 0x0980
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0988
    x"00",x"00",x"22",x"1C",x"22",x"22",x"22",x"22", -- 0x0990
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0998
    x"00",x"00",x"14",x"22",x"22",x"22",x"22",x"22", -- 0x09A0
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09A8
    x"00",x"00",x"1C",x"20",x"1C",x"22",x"1C",x"02", -- 0x09B0
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09B8
    x"00",x"00",x"04",x"0A",x"08",x"1C",x"08",x"0A", -- 0x09C0
    x"3C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09C8
    x"00",x"00",x"08",x"08",x"3E",x"08",x"08",x"00", -- 0x09D0
    x"3E",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09D8
    x"00",x"00",x"04",x"0A",x"04",x"00",x"00",x"00", -- 0x09E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09E8
    x"00",x"00",x"04",x"0A",x"08",x"1C",x"08",x"08", -- 0x09F0
    x"28",x"10",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A08
    x"00",x"00",x"08",x"08",x"08",x"08",x"08",x"00", -- 0x0A10
    x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A18
    x"00",x"00",x"14",x"14",x"14",x"00",x"00",x"00", -- 0x0A20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A28
    x"00",x"00",x"14",x"14",x"3E",x"14",x"3E",x"14", -- 0x0A30
    x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A38
    x"00",x"00",x"08",x"1E",x"28",x"1C",x"0A",x"3C", -- 0x0A40
    x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A48
    x"00",x"00",x"32",x"32",x"04",x"08",x"10",x"26", -- 0x0A50
    x"26",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A58
    x"00",x"00",x"10",x"28",x"28",x"10",x"2A",x"24", -- 0x0A60
    x"1A",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A68
    x"00",x"00",x"08",x"08",x"10",x"00",x"00",x"00", -- 0x0A70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A78
    x"00",x"00",x"08",x"10",x"20",x"20",x"20",x"10", -- 0x0A80
    x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A88
    x"00",x"00",x"08",x"04",x"02",x"02",x"02",x"04", -- 0x0A90
    x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A98
    x"00",x"00",x"00",x"08",x"2A",x"1C",x"1C",x"2A", -- 0x0AA0
    x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AA8
    x"00",x"00",x"00",x"08",x"08",x"3E",x"08",x"08", -- 0x0AB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08", -- 0x0AC0
    x"08",x"10",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AC8
    x"00",x"00",x"00",x"00",x"00",x"3E",x"00",x"00", -- 0x0AD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AE0
    x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AE8
    x"00",x"00",x"00",x"02",x"04",x"08",x"10",x"20", -- 0x0AF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AF8
    x"00",x"00",x"1C",x"22",x"26",x"2A",x"32",x"22", -- 0x0B00
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B08
    x"00",x"00",x"08",x"18",x"08",x"08",x"08",x"08", -- 0x0B10
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B18
    x"00",x"00",x"1C",x"22",x"02",x"1C",x"20",x"20", -- 0x0B20
    x"3E",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B28
    x"00",x"00",x"1C",x"22",x"02",x"04",x"02",x"22", -- 0x0B30
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B38
    x"00",x"00",x"04",x"0C",x"14",x"24",x"3E",x"04", -- 0x0B40
    x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B48
    x"00",x"00",x"3E",x"20",x"3C",x"02",x"02",x"02", -- 0x0B50
    x"3C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B58
    x"00",x"00",x"1C",x"20",x"20",x"3C",x"22",x"22", -- 0x0B60
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B68
    x"00",x"00",x"3E",x"02",x"04",x"08",x"10",x"20", -- 0x0B70
    x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B78
    x"00",x"00",x"1C",x"22",x"22",x"1C",x"22",x"22", -- 0x0B80
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B88
    x"00",x"00",x"1C",x"22",x"22",x"1E",x"02",x"02", -- 0x0B90
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B98
    x"00",x"00",x"00",x"00",x"08",x"00",x"00",x"08", -- 0x0BA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BA8
    x"00",x"00",x"00",x"00",x"08",x"00",x"00",x"08", -- 0x0BB0
    x"08",x"10",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BB8
    x"00",x"00",x"04",x"08",x"10",x"20",x"10",x"08", -- 0x0BC0
    x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BC8
    x"00",x"00",x"00",x"00",x"3E",x"00",x"3E",x"00", -- 0x0BD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BD8
    x"00",x"00",x"10",x"08",x"04",x"02",x"04",x"08", -- 0x0BE0
    x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BE8
    x"00",x"00",x"1C",x"22",x"02",x"04",x"08",x"00", -- 0x0BF0
    x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BF8
    x"00",x"00",x"1C",x"22",x"02",x"1A",x"2A",x"2A", -- 0x0C00
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C08
    x"00",x"00",x"08",x"14",x"22",x"22",x"3E",x"22", -- 0x0C10
    x"22",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C18
    x"00",x"00",x"3C",x"12",x"12",x"1C",x"12",x"12", -- 0x0C20
    x"3C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C28
    x"00",x"00",x"1C",x"22",x"20",x"20",x"20",x"22", -- 0x0C30
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C38
    x"00",x"00",x"3C",x"12",x"12",x"12",x"12",x"12", -- 0x0C40
    x"3C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C48
    x"00",x"00",x"3E",x"20",x"20",x"3C",x"20",x"20", -- 0x0C50
    x"3E",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C58
    x"00",x"00",x"3E",x"20",x"20",x"3C",x"20",x"20", -- 0x0C60
    x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C68
    x"00",x"00",x"1E",x"20",x"20",x"26",x"22",x"22", -- 0x0C70
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C78
    x"00",x"00",x"22",x"22",x"22",x"3E",x"22",x"22", -- 0x0C80
    x"22",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C88
    x"00",x"00",x"1C",x"08",x"08",x"08",x"08",x"08", -- 0x0C90
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C98
    x"00",x"00",x"02",x"02",x"02",x"02",x"22",x"22", -- 0x0CA0
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CA8
    x"00",x"00",x"22",x"24",x"28",x"30",x"28",x"24", -- 0x0CB0
    x"22",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CB8
    x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x0CC0
    x"3E",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CC8
    x"00",x"00",x"22",x"36",x"2A",x"2A",x"22",x"22", -- 0x0CD0
    x"22",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CD8
    x"00",x"00",x"22",x"32",x"2A",x"26",x"22",x"22", -- 0x0CE0
    x"22",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CE8
    x"00",x"00",x"1C",x"22",x"22",x"22",x"22",x"22", -- 0x0CF0
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CF8
    x"00",x"00",x"3C",x"22",x"22",x"3C",x"20",x"20", -- 0x0D00
    x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D08
    x"00",x"00",x"1C",x"22",x"22",x"22",x"2A",x"24", -- 0x0D10
    x"1A",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D18
    x"00",x"00",x"3C",x"22",x"22",x"3C",x"28",x"24", -- 0x0D20
    x"22",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D28
    x"00",x"00",x"1C",x"22",x"10",x"08",x"04",x"22", -- 0x0D30
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D38
    x"00",x"00",x"3E",x"08",x"08",x"08",x"08",x"08", -- 0x0D40
    x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D48
    x"00",x"00",x"22",x"22",x"22",x"22",x"22",x"22", -- 0x0D50
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D58
    x"00",x"00",x"22",x"22",x"22",x"14",x"14",x"08", -- 0x0D60
    x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D68
    x"00",x"00",x"22",x"22",x"22",x"2A",x"2A",x"36", -- 0x0D70
    x"22",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D78
    x"00",x"00",x"22",x"22",x"14",x"08",x"14",x"22", -- 0x0D80
    x"22",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D88
    x"00",x"00",x"22",x"22",x"14",x"08",x"08",x"08", -- 0x0D90
    x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D98
    x"00",x"00",x"3E",x"02",x"04",x"08",x"10",x"20", -- 0x0DA0
    x"3E",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DA8
    x"00",x"00",x"38",x"20",x"20",x"20",x"20",x"20", -- 0x0DB0
    x"38",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DB8
    x"00",x"00",x"20",x"20",x"10",x"08",x"04",x"02", -- 0x0DC0
    x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DC8
    x"00",x"00",x"0E",x"02",x"02",x"02",x"02",x"02", -- 0x0DD0
    x"0E",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DD8
    x"00",x"00",x"08",x"1C",x"2A",x"08",x"08",x"08", -- 0x0DE0
    x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DE8
    x"00",x"00",x"00",x"08",x"10",x"3E",x"10",x"08", -- 0x0DF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DF8
    x"00",x"00",x"08",x"14",x"22",x"00",x"00",x"00", -- 0x0E00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E08
    x"00",x"00",x"00",x"00",x"1C",x"02",x"1E",x"22", -- 0x0E10
    x"1E",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E18
    x"00",x"00",x"20",x"20",x"2C",x"32",x"22",x"32", -- 0x0E20
    x"2C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E28
    x"00",x"00",x"00",x"00",x"1C",x"22",x"20",x"22", -- 0x0E30
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E38
    x"00",x"00",x"02",x"02",x"1A",x"26",x"22",x"26", -- 0x0E40
    x"1A",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E48
    x"00",x"00",x"00",x"00",x"1C",x"22",x"3E",x"20", -- 0x0E50
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E58
    x"00",x"00",x"04",x"0A",x"08",x"1C",x"08",x"08", -- 0x0E60
    x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E68
    x"00",x"00",x"00",x"00",x"1A",x"26",x"26",x"1A", -- 0x0E70
    x"02",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E78
    x"00",x"00",x"20",x"20",x"2C",x"32",x"22",x"22", -- 0x0E80
    x"22",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E88
    x"00",x"00",x"00",x"08",x"00",x"18",x"08",x"08", -- 0x0E90
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E98
    x"00",x"00",x"00",x"02",x"00",x"02",x"02",x"02", -- 0x0EA0
    x"22",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EA8
    x"00",x"00",x"20",x"20",x"24",x"28",x"30",x"28", -- 0x0EB0
    x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EB8
    x"00",x"00",x"18",x"08",x"08",x"08",x"08",x"08", -- 0x0EC0
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EC8
    x"00",x"00",x"00",x"00",x"14",x"2A",x"2A",x"2A", -- 0x0ED0
    x"2A",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0ED8
    x"00",x"00",x"00",x"00",x"2C",x"32",x"22",x"22", -- 0x0EE0
    x"22",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EE8
    x"00",x"00",x"00",x"00",x"1C",x"22",x"22",x"22", -- 0x0EF0
    x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EF8
    x"00",x"00",x"00",x"00",x"2C",x"32",x"32",x"2C", -- 0x0F00
    x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F08
    x"00",x"00",x"00",x"00",x"1A",x"26",x"26",x"1A", -- 0x0F10
    x"02",x"02",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F18
    x"00",x"00",x"00",x"00",x"2C",x"32",x"20",x"20", -- 0x0F20
    x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F28
    x"00",x"00",x"00",x"00",x"1E",x"20",x"1C",x"02", -- 0x0F30
    x"3C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F38
    x"00",x"00",x"10",x"10",x"38",x"10",x"10",x"12", -- 0x0F40
    x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F48
    x"00",x"00",x"00",x"00",x"22",x"22",x"22",x"26", -- 0x0F50
    x"1A",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F58
    x"00",x"00",x"00",x"00",x"22",x"22",x"22",x"14", -- 0x0F60
    x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F68
    x"00",x"00",x"00",x"00",x"22",x"2A",x"2A",x"14", -- 0x0F70
    x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F78
    x"00",x"00",x"00",x"00",x"22",x"14",x"08",x"14", -- 0x0F80
    x"22",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F88
    x"00",x"00",x"00",x"00",x"22",x"22",x"22",x"1E", -- 0x0F90
    x"02",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F98
    x"00",x"00",x"00",x"00",x"3E",x"04",x"08",x"10", -- 0x0FA0
    x"3E",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FA8
    x"00",x"00",x"08",x"10",x"10",x"20",x"10",x"10", -- 0x0FB0
    x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FB8
    x"00",x"00",x"08",x"08",x"08",x"00",x"08",x"08", -- 0x0FC0
    x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FC8
    x"00",x"00",x"08",x"04",x"04",x"02",x"04",x"04", -- 0x0FD0
    x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FD8
    x"00",x"00",x"10",x"2A",x"04",x"00",x"00",x"00", -- 0x0FE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FF0
    x"3E",x"00",x"00",x"00",x"00",x"00",x"00",x"00"  -- 0x0FF8
  );

begin

  p_rom_wr:		process
				begin
				wait until rising_edge(WR_CLK);
					if WE = '1' then
						RAM(to_integer(unsigned(ADDR_W))) <= DATA_W;
					end if;
				end process;

  p_rom_rd:		process
				begin
				wait until rising_edge(RD_CLK);
					DATA_R <= RAM(to_integer(unsigned(ADDR_R)));
				end process;

end RTL;
