 #            ����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ����  �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  �2NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  	s�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  �PNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  P�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  �_NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  
&�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  6�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  �,NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  �aNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  @�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  �nNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  �NNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  c�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� sMNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� &NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
PBNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� @|NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ژNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 6 NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� csNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� /NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� dNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ZNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� a8NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� B7NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 4kNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
˞NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ۠NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ADNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� R	NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� qNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� '&NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� a�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� q�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	�yNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �%NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� b�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �vNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 4�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� B�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
�*NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 7�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� $�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �HNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� Q�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �GNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� 0�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	�TNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 3�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� F�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �[NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� e�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �9NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� f�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� u�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �eNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� V�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �6NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �jNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� FINNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� VwNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� E:NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 0NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� eFNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� iNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� $NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  +NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� vNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� ݕNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ͫNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	T<NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� "`NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� w3NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
oNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� QNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� gNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 2^NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� DNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� �!NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	"�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� T�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �RNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �}NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �rNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �.NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
w�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� g�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �LNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �CNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �cNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� D�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 2�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� o�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	�fNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �:NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� |�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �iNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� *�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� \�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
�5NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� )�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� :�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �WNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� O�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �XNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ����	 	{NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����	 ENNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����	 	��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����	 ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����	 
NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����	 'NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����	 ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����	 \(NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����	 *tNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����	 
ՁNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����	 ſNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����	 _[NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����	 LNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����	 ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����	 oNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����	 99NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����	 �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����	 ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ����
 ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����
 ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����
 	NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����
 mRNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����
 ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����
 ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����
 8NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����
 ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����
 ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����
 
N]NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����
 ^cNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����
 ćNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����
 ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����
 (?NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����
 ��NNNNNNNNNNNNNNNNNNNNNN            ������������������������������������������������������������������������������������������������������������������������������������������������������������������& V�1.0 & 
� 80 & � &' LS$�"  " &6 (� &HFFD9,0 &u 2� SUNDAY,MONDAY,TUESDAY,WEDNESDAY,THURSDAY,FRIDAY,SATURDAY &� <� JAN,FEB,MAR,APR,MAY,JUN,JUL,AUG,SEPT,OCT,NOV,DEC &� FY���(&HFFC0)�100���(&HFFC1) &� PMN���(&HFFC2) &� ZDM���(&HFFC3) ' dDW���(&HFFC4) ' nHR���(&HFFC5) '& xMI���(&HFFC6) '7 �S���(&HFFC7) 'B ��� 160 'M ��� 250 '] ��:� A�1 � 7 'f �� F$ 'y �� A�DW � D$�F$ '� �� A '� Ȁ A�1 � 12 '� ҍ F$ '� ܅ A�MN � N$�F$ '� � '� � '� �� '�� HR � 10 � HR$�"0"���(��(HR),1) :� HR$���(��(HR),2) (0� MI � 10 � MI$�"0"���(��(MI),1) :� MI$���(��(MI),2) (d� S � 10 � S$�"0"���(��(S),1) :� S$���(��(S),2) (w"� LS$�S$ � 310 (�,�� 340 (�6LS$�S$ (�J�� 70 (�T� 0,0 (�^� "Today is: ";D$ (�h� N$;" ";DM;" ";Y (�r� HR$;" : ";MI$;" : ";S$ (�|�   ),2) (0� M����������NNNNNNNNNNNNNNNNNNNNNNNN        ����
 0NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �-NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	m�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �`NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �ONNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� N�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �@NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
8�NNNNNNNNNNNNNNNNNNNNNN            ������������������������������������������������������������&	 I�0 & V�1.2 & 
� D(16) &7 � @192,"         "; &O � @128,"ID VER=";V; &Z (�� 340 &� -� DB�1 � � " *** DEBUG MODE ***" :� � "" &� 2� D(10) �� 10 � 330 &� <V$�" 20" &� F� X�1 � 9 &� PV$�V$���(D(X)) &� Z� X�6 � V$�V$�"-" &� _� X�2 � V$�V$�"." ' `� X�4 � V$�V$�"." ' d� X '2 n� "MISTER COCO3 V:";V$ 'B xLSB�0:MSB�0 '_ �� (D(12) � 1) �0 � LSB�1 '| �� (D(12) � 2) �0 � MSB�1 '� �M$�"" '� �� LSB � 0 � MSB � 1 � M$�"64MB" '� �� LSB�1 � MSB�0 � M$�"32MB" '� �� LSB�1 � MSB�1 � M$�"128MB" ( �� "MISTER MEMORY = ";M$;" SDRAM..." (' ȇ "BUILD CFG:"; (: Ҁ X�7 � 0 � �1 (e ܅ (D(11) � (2�X))�0 � F(X)�1 :� F(X)�0 (k � (v �F$�"(" (� �� X�1 � 8 (�� F(X�1)�1 � F$�F$���(��(X),1) :� F$�F$�" " (�� (�F$�F$�")" (�"� F$;" "; (�,� X�13 � 14 (�6� "$";��(D(X));" "; )@� )C� DB�1 � 330 )CE� @128,"                               "; )RF� @256,""; )eJ� I�1 � � :� � )tT� X�1 � 16 )�^D(X) � ��(&HFFEF) )�r� )�s� D(10) �128 � DB�1 )�tD(10) � D(10) � 15 )�|� )�� RUN 1000 TO DEBUG )��I�1:�:�� 5   ";��(D(X));" "; ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ^�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �qNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �QNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN        �c& V�1.1 & 
� &HFFD9,0 &@ � 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0 &v � 126,129,165,129,189,153,129,126,0,0,0,0,0,0,0,0 &� (� 126,255,219,255,195,231,255,126,0,0,0,0,0,0,0,0 &� 2� 108,254,254,254,124,56,16,0,0,0,0,0,0,0,0,0 ' <� 16,56,124,254,124,56,16,0,0,0,0,0,0,0,0,0 'A F� 56,124,56,254,254,124,56,124,0,0,0,0,0,0,0,0 's P� 16,16,56,124,254,124,56,124,0,0,0,0,0,0,0,0 '� Z� 0,0,24,60,60,24,0,0,0,0,0,0,0,0,0,0 '� d� 255,255,231,195,195,231,255,255,0,0,0,0,0,0,0,0 ( n� 0,60,102,66,66,102,60,0,0,0,0,0,0,0,0,0 (7 x� 255,195,153,189,189,153,195,255,0,0,0,0,0,0,0,0 (i �� 15,7,15,125,204,204,204,120,0,0,0,0,0,0,0,0 (� �� 60,102,102,102,60,24,126,24,0,0,0,0,0,0,0,0 (� �� 63,51,63,48,48,112,240,224,0,0,0,0,0,0,0,0 (� �� 127,99,127,99,99,103,230,192,0,0,0,0,0,0,0,0 )1 �� 153,90,60,231,231,60,90,153,0,0,0,0,0,0,0,0 )e �� 128,224,248,254,248,224,128,0,0,0,0,0,0,0,0,0 )� �� 2,14,62,254,62,14,2,0,0,0,0,0,0,0,0,0 )� Ȇ 24,60,126,24,24,126,60,24,0,0,0,0,0,0,0,0 )� ҆ 102,102,102,102,102,0,102,0,0,0,0,0,0,0,0,0 *$ ܆ 127,219,219,123,27,27,27,0,0,0,0,0,0,0,0,0 *W � 60,102,56,108,108,56,204,120,0,0,0,0,0,0,0,0 *� �� 0,0,0,0,126,126,126,0,0,0,0,0,0,0,0,0 *� �� 24,60,126,24,126,60,24,255,0,0,0,0,0,0,0,0 *�� 24,60,126,24,24,24,24,0,0,0,0,0,0,0,0,0 +� 24,24,24,24,126,60,24,0,0,0,0,0,0,0,0,0 +<� 0,24,12,254,12,24,0,0,0,0,0,0,0,0,0,0 +h"� 0,48,96,254,96,48,0,0,0,0,0,0,0,0,0,0 +�,� 0,0,192,192,192,254,0,0,0,0,0,0,0,0,0,0 +�6� 0,36,102,255,102,36,0,0,0,0,0,0,0,0,0,0 +�@� 0,24,60,126,255,255,0,0,0,0,0,0,0,0,0,0 , J� 0,255,255,126,60,24,0,0,0,0,0,0,0,0,0,0 ,FT� 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0 ,t^� 48,120,120,48,48,0,48,0,0,0,0,0,0,0,0,0 ,�h� 108,108,108,0,0,0,0,0,0,0,0,0,0,0,0,0 ,�r� 108,108,254,108,254,108,108,0,0,0,0,0,0,0,0,0 -|� 48,124,192,120,12,248,48,0,0,0,0,0,0,0,0,0 -5�� 0,198,204,24,48,102,198,0,0,0,0,0,0,0,0,0 -g�� 56,108,56,118,220,204,118,0,0,0,0,0,0,0,0,0 -��� 96,96,192,0,0,0,0,0,0,0,0,0,0,0,0,0 -��� 24,48,96,96,96,48,24,0,0,0,0,0,0,0,0,0 -��� 96,48,24,24,24,48,96,0,0,0,0,0,0,0,0,0 .�� 0,102,60,255,60,102,0,0,0,0,0,0,0,0,0,0 .E 0,48,48,252,48,48,0,0,0,0,0,0,0,0,0,0 .n̆ 0,0,0,0,0,48,48,96,0,0,0,0,0,0,0,0 .�ֆ 0,0,0,252,0,0,0,0,0,0,0,0,0,0,0,0 .��� 0,0,0,0,0,48,48,0,0,0,0,0,0,0,0,0 .�� 6,12,24,48,96,192,128,0,0,0,0,0,0,0,0,0 / � 124,198,206,���� �MNNNNNNNNNNNNNNNNNNNNNN            �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������"#���������������NNNNNNNNNNNNNNNNNN                                                                                                                                                                                            AUTO    BAS    �                IBMFONT BAS  ! f                TESTRTC BAS   �                ������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �mNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �1NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
i�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� y�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �SNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �\NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �|NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� Z�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ,�NNNNNNNNNNNNNNNNNNNNNN            ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������222,246,230,124,0,0,0,0,0,0,0,0,0 /N�� 48,112,48,48,48,48,48,0,0,0,0,0,0,0,0,0 /� 120,204,12,56,96,192,252,0,0,0,0,0,0,0,0,0 /�� 120,204,12,56,12,204,120,0,0,0,0,0,0,0,0,0 /�� 28,60,108,204,254,12,12,0,0,0,0,0,0,0,0,0 0&� 252,192,248,12,12,204,120,0,0,0,0,0,0,0,0,0 0D0� 56,96,192,248,204,204,120,0,0,0,0,0,0,0,0,0 0r:� 252,12,12,24,48,48,48,0,0,0,0,0,0,0,0,0 0�D� 120,204,204,120,204,204,120,0,0,0,0,0,0,0,0,0 0�N� 120,204,204,124,12,24,112,0,0,0,0,0,0,0,0,0 1X� 0,48,48,0,0,48,48,0,0,0,0,0,0,0,0,0 1-b� 0,48,48,0,0,48,48,96,0,0,0,0,0,0,0,0 1[l� 24,48,96,192,96,48,24,0,0,0,0,0,0,0,0,0 1�v� 0,0,252,0,0,252,0,0,0,0,0,0,0,0,0,0 1��� 96,48,24,12,24,48,96,0,0,0,0,0,0,0,0,0 1��� 120,204,12,24,48,0,48,0,0,0,0,0,0,0,0,0 2�� 124,198,222,222,222,192,120,0,0,0,0,0,0,0,0,0 2F�� 24,60,102,102,126,102,102,0,0,0,0,0,0,0,0,0 2z�� 124,102,102,124,102,102,124,0,0,0,0,0,0,0,0,0 2��� 60,102,192,192,192,102,60,0,0,0,0,0,0,0,0,0 2��� 120,108,102,102,102,108,120,0,0,0,0,0,0,0,0,0 3Ɔ 126,96,96,120,96,96,126,0,0,0,0,0,0,0,0,0 3?І 126,96,96,120,96,96,96,0,0,0,0,0,0,0,0,0 3qچ 60,102,192,192,206,102,62,0,0,0,0,0,0,0,0,0 3�� 102,102,102,126,102,102,102,0,0,0,0,0,0,0,0,0 3�� 24,24,24,24,24,24,24,0,0,0,0,0,0,0,0,0 3��� 6,6,6,6,102,102,60,0,0,0,0,0,0,0,0,0 41� 102,102,108,120,108,102,102,0,0,0,0,0,0,0,0,0 4_� 96,96,96,96,96,96,126,0,0,0,0,0,0,0,0,0 4�� 198,238,254,254,214,198,198,0,0,0,0,0,0,0,0,0 4� � 198,230,246,222,206,198,198,0,0,0,0,0,0,0,0,0 4�*� 60,102,102,102,102,102,60,0,0,0,0,0,0,0,0,0 5*4� 124,102,102,124,96,96,96,0,0,0,0,0,0,0,0,0 5[>� 60,102,102,102,110,60,14,0,0,0,0,0,0,0,0,0 5�H� 124,102,102,124,108,102,102,0,0,0,0,0,0,0,0,0 5�R� 60,102,112,56,14,102,60,0,0,0,0,0,0,0,0,0 5�\� 126,24,24,24,24,24,24,0,0,0,0,0,0,0,0,0 6 f� 102,102,102,102,102,102,62,0,0,0,0,0,0,0,0,0 6Rp� 102,102,102,102,102,60,24,0,0,0,0,0,0,0,0,0 6�z� 198,198,198,214,254,238,198,0,0,0,0,0,0,0,0,0 6��� 102,102,60,24,60,102,102,0,0,0,0,0,0,0,0,0 6��� 102,102,102,60,24,24,24,0,0,0,0,0,0,0,0,0 7�� 254,6,12,24,48,96,254,0,0,0,0,0,0,0,0,0 7D�� 120,96,96,96,96,96,120,0,0,0,0,0,0,0,0,0 7p�� 192,96,48,24,12,6,2,0,0,0,0,0,0,0,0,0 7��� 120,24,24,24,24,24,120,0,0,0,0,0,0,0,0,0 7��� 16,56,108,198,0,0,0,0,0,0,0,0,0,0,0,0 7�ʆ 0,0,0,0,0,0,0,255,0,0,0,0,0,0,0,0 8Ԇ 48,48,24,0,0,0,0,0,0,0,0,0,0,0,0,0 8Gކ 0,0,60,6,62,102,58,0,0,0,0,0,0,0,0,0 8w� 96,96,96,124,102,102,92,0,0,0,0,0,0,0,0,0 8�� 0,0,60,102,96,102,60,0,0,0,0,0,0,0,0,0 8��� 6,6,6,62,102,102,58,0,0,0,0,0,0,0,0,0 8�� 0,0,60,102,126,96,60,0,0,0,0,0,0,0,0,0 9+� 28,54,48,120,48,48,48,0,0,0,0,0,0,0,0,0 9X� 0,0,58,102,102,62,6,60,0,0,0,0,0,0,0,0 9�$� 96,96,108,118,102,102,102,0,0,0,0,0,0,0,0,0 9�.� 24,0,24,24,24,24,24,0,0,0,0,0,0,0,0,0 9�8� 12,0,12,12,12,204,204,120,0,0,0,0,0,0,0,0 :B� 96,96,102,108,120,108,102,0,0,0,0,0,0,0,0,0 :EL� 24,24,24,24,24,24,24,0,0,0,0,0,0,0,0,0 :uV� 0,0,198,238,254,214,198,0,0,0,0,0,0,0,0,0 :�`� 0,0,124,102,102,102,102,0,0,0,0,0,0,0,0,0 :�j� 0,0,60,102,102,102,60,0,0,0,0,0,0,0,0,0 ;t� 0,0,92,102,102,124,96,96,0,0,0,0,0,0,0,0 ;.~� 0,0,58,102,102,62,6,6,0,0,0,0,0,0,0,0 ;Z�� 0,0,92,118,96,96,96,0,0,0,0,0,0,0,0,0 ;��� 0,0,62,96,60,6,124,0,0,0,0,0,0,0,0,0 ;��� 48,48,124,48,48,52,24,0,0,0,0,0,0,0,0,0 ;��� 0,0,102,102,102,102,58,0,0,0,0,0,0,0,0,0 <�� 0,0,102,102,102,60,24,0,0,0,0,0,0,0,0,0 <@�� 0,0,198,214,254,254,108,0,0,0,0,0,0,0,0,0 <oĆ 0,0,198,108,58,108,198,0,0,0,0,0,0,0,0,0 <�Ά 0,0,102,102,102,62,6,60,0,0,0,0,0,0,0,0 <�؆ 0,0,126,12,24,48,126,0,0,0,0,0,0,0,0,0 <�� 28,48,48,224,48,48,28,0,0,0,0,0,0,0,0,0 =$� 24,24,24,0,24,24,24,0,0,0,0,0,0,0,0,0 =S�� 224,48,48,28,48,48,224,0,0,0,0,0,0,0,0,0 =} � 118,220,0,0,0,0,0,0,0,0,0,0,0,0,0,0 =�
� 0,16,56,108,198,198,254,0,0,0,0,0,0,0,0,0 =�� &HFFF0,&H5A =�� A � 0 � 2047 =�(� B =�2� &HFFF1,B =�<� A > F� &HFFF0,0 >P�80 >Z� >dB�0 >6n� A � &H6C000 � A � 511 � 4 >@x� A,B >J�B�B�1 >R�� A >\�� 1,8 >b��   ,0,0,0,0,0,0,0,0,0,0,0,0 =�
� 0,16,56,108,198,198,254,0,0,0,0,0,0,0,0,0 =�� &HFFF0,&H5A =�� A � 0 � 2047 =�(� B =�2� &HFFF1,B =�<� A > F� &HFFF0,������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� yNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ,ANNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ZNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� XVNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� HhNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� [%NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� .
NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� {YNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� vNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ;NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� >4NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� hNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� .�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� >�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	�KNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� -�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� X�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �DNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� {�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �&NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� x�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� k�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �zNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� H�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �)NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �uNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	hNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ^NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� KNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ¤NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
=QNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� -oNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� [3NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� `NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� x<NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �!NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� h�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �lNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �CNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� =�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �LNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
K�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� [�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �?NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �rNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� -�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �}NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �]NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� x�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	�jNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �6NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� z�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �eNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� Y�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� /�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
�9NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� Z�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� I�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �[NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� j�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� <�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �TNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� zwNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� jINNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� yNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� +NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� /$NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� YxNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ,WNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ?NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� J5NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� +ZNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ;dNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ԯNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ()NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ]NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ~	NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� UNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� }zNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� n7NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� M8NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� đNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� ]�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� M�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	�GNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ^�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� +�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �HNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ~�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �*NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �vNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ;�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� m�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �%NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �yNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� �2NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	O�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 9�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �ANNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �nNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� l�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �aNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �=NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �_NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� |�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �PNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �pNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� )�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� _�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	9/NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� OsNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
l|NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� |BNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� _MNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� )NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� dhNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� tVNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� gNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 4NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 1;NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� GgNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 2HNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� !NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� T*NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	�uNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �)NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� d�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �zNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� G�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 1�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
�&NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� D�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� W�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �DNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� t�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� "�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �KNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� � NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �>NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	 �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� v�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �sNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �\NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� #�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �SNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
U�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� E�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� � NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �mNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 3�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �bNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �BNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� f�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	vNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  ANNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� UNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ܻNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
#NNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 3pNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� E,NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� f#NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	'0NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� QlNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ?NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
rcNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� b]NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ARNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 7NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� �-NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	Q�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� '�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �^NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �qNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� r�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �~NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �"NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �@NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� b�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �ONNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �oNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 7�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� A�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� C�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� S�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	�XNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� @�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 5�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �WNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� `�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �5NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �iNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� %�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� s�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �:NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� �fNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ���� 5ENNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� %{NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 	��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ʰNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 66NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� CNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� `NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� JNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� 
�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ceNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� p(NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� S'NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ڎNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ���� ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ����  �BNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  �|NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  	D�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  2�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  �1NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  g�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  �MNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  
�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  �bNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  �/NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  w�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  � NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  � NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  "�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����  T�NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ����! ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����! ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����! 	2_NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����! DNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����! ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����! ͪNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����! PNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����! �NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����! ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����! 
gNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����! w2NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����! ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����! ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����! nNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����! ݔNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����! ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����! T=NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����! "aNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN����O����E����;���ߍ1���Ց'�y�˕�                                                                                            NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN        ����"  *NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����" 0NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����" 	��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����" ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����" #YNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����" VvNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����" ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����" uyNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����" %NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����" 
��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����" ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����" v
NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����" eGNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����" ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����" FHNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����" hNNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����" ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNN        ����" ��NNNNNNNNNNNNNNNNNNNNNN            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN